`include "svmock_pkg.sv"

package ut_pkg;
  import svmock_pkg::*;

  `include "call.sv"
  `include "mock_call.sv"
endpackage
