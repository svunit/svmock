class call;

endclass
