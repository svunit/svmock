class mock_call extends call;

endclass
