module test(
  input            clk,
  input            rst_n,

  input            bit_i,
  input      [7:0] byte_i,
  output reg       bit_o,
  output reg [7:0] byte_o
);

endmodule
