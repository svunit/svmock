class bedrock;
  flintstones f = new();

  function void yabba_dabda_do(string wilma [int]);
    f.dino();
    f.bam_bam(f.pebbles(wilma.num(), wilma));
  endfunction
endclass
