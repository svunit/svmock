package svmock_pkg;
endpackage
