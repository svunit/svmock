class flintstones;
  function new(); endfunction

  function void dino();
    // all the code for dino
  endfunction

  function int pebbles(int fred, string wilma [int]);
    return 12;
  endfunction

  function void bam_bam(int barney);
    // nothing to do
  endfunction
endclass
