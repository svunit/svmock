`define SVMOCK_VOIDFUNCTION0(NAME) \
__mocker0 #() __``NAME = new("NAME", __mockers); \
function NAME(); \
  __``NAME.Called(); \
  super.NAME(); \
endfunction

`define SVMOCK_FUNCTION0(NAME, RETURN) \
__mocker0 #() __``NAME = new("NAME", __mockers); \
function RETURN NAME(); \
  __``NAME.Called(); \
  return super.NAME(); \
endfunction

`define SVMOCK_VOIDFUNCTION1(NAME,TYPE0,ARG0) \
__mocker1 #(TYPE0) __``NAME = new("NAME", __mockers); \
function NAME(TYPE0 ARG0); \
  __``NAME.Called(ARG0); \
  super.NAME(ARG0); \
endfunction

`define SVMOCK_FUNCTION1(NAME, RETURN,TYPE0,ARG0) \
__mocker1 #(TYPE0) __``NAME = new("NAME", __mockers); \
function RETURN NAME(TYPE0 ARG0); \
  __``NAME.Called(ARG0); \
  return super.NAME(ARG0); \
endfunction

`define SVMOCK_VOIDFUNCTION2(NAME,TYPE0,ARG0,TYPE1,ARG1) \
__mocker2 #(TYPE0, TYPE1) __``NAME = new("NAME", __mockers); \
function NAME(TYPE0 ARG0, TYPE1 ARG1); \
  __``NAME.Called(ARG0,ARG1); \
  super.NAME(ARG0,ARG1); \
endfunction

`define SVMOCK_FUNCTION2(NAME, RETURN,TYPE0,ARG0,TYPE1,ARG1) \
__mocker2 #(TYPE0, TYPE1) __``NAME = new("NAME", __mockers); \
function RETURN NAME(TYPE0 ARG0, TYPE1 ARG1); \
  __``NAME.Called(ARG0,ARG1); \
  return super.NAME(ARG0,ARG1); \
endfunction

`define SVMOCK_VOIDFUNCTION3(NAME,TYPE0,ARG0,TYPE1,ARG1,TYPE2,ARG2) \
__mocker3 #(TYPE0, TYPE1, TYPE2) __``NAME = new("NAME", __mockers); \
function NAME(TYPE0 ARG0, TYPE1 ARG1, TYPE2 ARG2); \
  __``NAME.Called(ARG0,ARG1,ARG2); \
  super.NAME(ARG0,ARG1,ARG2); \
endfunction

`define SVMOCK_FUNCTION3(NAME, RETURN,TYPE0,ARG0,TYPE1,ARG1,TYPE2,ARG2) \
__mocker3 #(TYPE0, TYPE1, TYPE2) __``NAME = new("NAME", __mockers); \
function RETURN NAME(TYPE0 ARG0, TYPE1 ARG1, TYPE2 ARG2); \
  __``NAME.Called(ARG0,ARG1,ARG2); \
  return super.NAME(ARG0,ARG1,ARG2); \
endfunction

`define SVMOCK_VOIDFUNCTION4(NAME,TYPE0,ARG0,TYPE1,ARG1,TYPE2,ARG2,TYPE3,ARG3) \
__mocker4 #(TYPE0, TYPE1, TYPE2, TYPE3) __``NAME = new("NAME", __mockers); \
function NAME(TYPE0 ARG0, TYPE1 ARG1, TYPE2 ARG2, TYPE3 ARG3); \
  __``NAME.Called(ARG0,ARG1,ARG2,ARG3); \
  super.NAME(ARG0,ARG1,ARG2,ARG3); \
endfunction

`define SVMOCK_FUNCTION4(NAME, RETURN,TYPE0,ARG0,TYPE1,ARG1,TYPE2,ARG2,TYPE3,ARG3) \
__mocker4 #(TYPE0, TYPE1, TYPE2, TYPE3) __``NAME = new("NAME", __mockers); \
function RETURN NAME(TYPE0 ARG0, TYPE1 ARG1, TYPE2 ARG2, TYPE3 ARG3); \
  __``NAME.Called(ARG0,ARG1,ARG2,ARG3); \
  return super.NAME(ARG0,ARG1,ARG2,ARG3); \
endfunction

`define SVMOCK_VOIDFUNCTION5(NAME,TYPE0,ARG0,TYPE1,ARG1,TYPE2,ARG2,TYPE3,ARG3,TYPE4,ARG4) \
__mocker5 #(TYPE0, TYPE1, TYPE2, TYPE3, TYPE4) __``NAME = new("NAME", __mockers); \
function NAME(TYPE0 ARG0, TYPE1 ARG1, TYPE2 ARG2, TYPE3 ARG3, TYPE4 ARG4); \
  __``NAME.Called(ARG0,ARG1,ARG2,ARG3,ARG4); \
  super.NAME(ARG0,ARG1,ARG2,ARG3,ARG4); \
endfunction

`define SVMOCK_FUNCTION5(NAME, RETURN,TYPE0,ARG0,TYPE1,ARG1,TYPE2,ARG2,TYPE3,ARG3,TYPE4,ARG4) \
__mocker5 #(TYPE0, TYPE1, TYPE2, TYPE3, TYPE4) __``NAME = new("NAME", __mockers); \
function RETURN NAME(TYPE0 ARG0, TYPE1 ARG1, TYPE2 ARG2, TYPE3 ARG3, TYPE4 ARG4); \
  __``NAME.Called(ARG0,ARG1,ARG2,ARG3,ARG4); \
  return super.NAME(ARG0,ARG1,ARG2,ARG3,ARG4); \
endfunction

`define SVMOCK_VOIDFUNCTION6(NAME,TYPE0,ARG0,TYPE1,ARG1,TYPE2,ARG2,TYPE3,ARG3,TYPE4,ARG4,TYPE5,ARG5) \
__mocker6 #(TYPE0, TYPE1, TYPE2, TYPE3, TYPE4, TYPE5) __``NAME = new("NAME", __mockers); \
function NAME(TYPE0 ARG0, TYPE1 ARG1, TYPE2 ARG2, TYPE3 ARG3, TYPE4 ARG4, TYPE5 ARG5); \
  __``NAME.Called(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5); \
  super.NAME(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5); \
endfunction

`define SVMOCK_FUNCTION6(NAME, RETURN,TYPE0,ARG0,TYPE1,ARG1,TYPE2,ARG2,TYPE3,ARG3,TYPE4,ARG4,TYPE5,ARG5) \
__mocker6 #(TYPE0, TYPE1, TYPE2, TYPE3, TYPE4, TYPE5) __``NAME = new("NAME", __mockers); \
function RETURN NAME(TYPE0 ARG0, TYPE1 ARG1, TYPE2 ARG2, TYPE3 ARG3, TYPE4 ARG4, TYPE5 ARG5); \
  __``NAME.Called(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5); \
  return super.NAME(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5); \
endfunction

`define SVMOCK_VOIDFUNCTION7(NAME,TYPE0,ARG0,TYPE1,ARG1,TYPE2,ARG2,TYPE3,ARG3,TYPE4,ARG4,TYPE5,ARG5,TYPE6,ARG6) \
__mocker7 #(TYPE0, TYPE1, TYPE2, TYPE3, TYPE4, TYPE5, TYPE6) __``NAME = new("NAME", __mockers); \
function NAME(TYPE0 ARG0, TYPE1 ARG1, TYPE2 ARG2, TYPE3 ARG3, TYPE4 ARG4, TYPE5 ARG5, TYPE6 ARG6); \
  __``NAME.Called(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5,ARG6); \
  super.NAME(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5,ARG6); \
endfunction

`define SVMOCK_FUNCTION7(NAME, RETURN,TYPE0,ARG0,TYPE1,ARG1,TYPE2,ARG2,TYPE3,ARG3,TYPE4,ARG4,TYPE5,ARG5,TYPE6,ARG6) \
__mocker7 #(TYPE0, TYPE1, TYPE2, TYPE3, TYPE4, TYPE5, TYPE6) __``NAME = new("NAME", __mockers); \
function RETURN NAME(TYPE0 ARG0, TYPE1 ARG1, TYPE2 ARG2, TYPE3 ARG3, TYPE4 ARG4, TYPE5 ARG5, TYPE6 ARG6); \
  __``NAME.Called(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5,ARG6); \
  return super.NAME(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5,ARG6); \
endfunction

`define SVMOCK_VOIDFUNCTION8(NAME,TYPE0,ARG0,TYPE1,ARG1,TYPE2,ARG2,TYPE3,ARG3,TYPE4,ARG4,TYPE5,ARG5,TYPE6,ARG6,TYPE7,ARG7) \
__mocker8 #(TYPE0, TYPE1, TYPE2, TYPE3, TYPE4, TYPE5, TYPE6, TYPE7) __``NAME = new("NAME", __mockers); \
function NAME(TYPE0 ARG0, TYPE1 ARG1, TYPE2 ARG2, TYPE3 ARG3, TYPE4 ARG4, TYPE5 ARG5, TYPE6 ARG6, TYPE7 ARG7); \
  __``NAME.Called(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5,ARG6,ARG7); \
  super.NAME(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5,ARG6,ARG7); \
endfunction

`define SVMOCK_FUNCTION8(NAME, RETURN,TYPE0,ARG0,TYPE1,ARG1,TYPE2,ARG2,TYPE3,ARG3,TYPE4,ARG4,TYPE5,ARG5,TYPE6,ARG6,TYPE7,ARG7) \
__mocker8 #(TYPE0, TYPE1, TYPE2, TYPE3, TYPE4, TYPE5, TYPE6, TYPE7) __``NAME = new("NAME", __mockers); \
function RETURN NAME(TYPE0 ARG0, TYPE1 ARG1, TYPE2 ARG2, TYPE3 ARG3, TYPE4 ARG4, TYPE5 ARG5, TYPE6 ARG6, TYPE7 ARG7); \
  __``NAME.Called(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5,ARG6,ARG7); \
  return super.NAME(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5,ARG6,ARG7); \
endfunction

`define SVMOCK_VOIDFUNCTION9(NAME,TYPE0,ARG0,TYPE1,ARG1,TYPE2,ARG2,TYPE3,ARG3,TYPE4,ARG4,TYPE5,ARG5,TYPE6,ARG6,TYPE7,ARG7,TYPE8,ARG8) \
__mocker9 #(TYPE0, TYPE1, TYPE2, TYPE3, TYPE4, TYPE5, TYPE6, TYPE7, TYPE8) __``NAME = new("NAME", __mockers); \
function NAME(TYPE0 ARG0, TYPE1 ARG1, TYPE2 ARG2, TYPE3 ARG3, TYPE4 ARG4, TYPE5 ARG5, TYPE6 ARG6, TYPE7 ARG7, TYPE8 ARG8); \
  __``NAME.Called(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5,ARG6,ARG7,ARG8); \
  super.NAME(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5,ARG6,ARG7,ARG8); \
endfunction

`define SVMOCK_FUNCTION9(NAME, RETURN,TYPE0,ARG0,TYPE1,ARG1,TYPE2,ARG2,TYPE3,ARG3,TYPE4,ARG4,TYPE5,ARG5,TYPE6,ARG6,TYPE7,ARG7,TYPE8,ARG8) \
__mocker9 #(TYPE0, TYPE1, TYPE2, TYPE3, TYPE4, TYPE5, TYPE6, TYPE7, TYPE8) __``NAME = new("NAME", __mockers); \
function RETURN NAME(TYPE0 ARG0, TYPE1 ARG1, TYPE2 ARG2, TYPE3 ARG3, TYPE4 ARG4, TYPE5 ARG5, TYPE6 ARG6, TYPE7 ARG7, TYPE8 ARG8); \
  __``NAME.Called(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5,ARG6,ARG7,ARG8); \
  return super.NAME(ARG0,ARG1,ARG2,ARG3,ARG4,ARG5,ARG6,ARG7,ARG8); \
endfunction

