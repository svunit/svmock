package bedrock_pkg;
  `include "flintstones.sv"
  `include "bedrock.sv"
endpackage
