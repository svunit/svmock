`SVMOCK(mock_flintstones, flintstones)
  `SVMOCK_VFUNC0(dino)
  `SVMOCK_FUNC2(pebbles, int, int, fred, , string, wilma, [int])
  `SVMOCK_VFUNC1(bam_bam, int, barney, )
`SVMOCK_END
