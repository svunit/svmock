class apb_item extends uvm_sequence_item;
endclass
