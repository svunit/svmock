`SVMOCK(mock_flintstones, flintstones)
  `SVMOCK_VOIDFUNCTION0(dino)
  `SVMOCK_FUNCTION2(pebbles, int, int, fred, , string, wilma, [int])
  `SVMOCK_VOIDFUNCTION1(bam_bam, int, barney, )
`SVMOCK_END
